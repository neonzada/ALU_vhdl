library verilog;
use verilog.vl_types.all;
entity ULAcompleta_vlg_vec_tst is
end ULAcompleta_vlg_vec_tst;
